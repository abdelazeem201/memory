# 
# LEF OUT 
# User Name : rimah 
# Date : Tue Sep 28 12:54:50 2010
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SRAM16x64
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 154.59 BY 160.505 ;
  SYMMETRY X Y R90 ;

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 35.135 0.16 35.295 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 35.135 0.16 35.295 ;
    END
  END WEB2

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.43 34.065 154.59 34.225 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.43 34.065 154.59 34.225 ;
    END
  END WEB1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 129.25 0 133.25 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.455 0 145.455 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.495 0 67.495 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.41 0 78.41 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.385 0 100.385 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.305 0 111.305 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.95 0 45.95 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.41 0 11.41 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.45 0 23.45 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.95 156.505 45.95 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.495 156.505 67.495 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.41 156.505 78.41 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.385 156.505 100.385 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.305 156.505 111.305 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.25 156.505 133.25 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.455 156.505 145.455 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.45 156.505 23.45 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.41 156.505 11.41 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.45 0 23.45 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.305 0 111.305 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.41 0 11.41 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.95 0 45.95 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.25 0 133.25 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.495 0 67.495 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.385 0 100.385 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.41 0 78.41 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.455 0 145.455 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.95 156.505 45.95 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.495 156.505 67.495 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.41 156.505 78.41 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.385 156.505 100.385 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.305 156.505 111.305 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.25 156.505 133.25 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.455 156.505 145.455 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.45 156.505 23.45 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.41 156.505 11.41 160.505 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 112.615 0 116.615 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.26 0 51.26 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.56 0 138.56 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.72 0 83.72 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.765 0 150.765 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.46 0 5.46 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.76 0 28.76 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.695 0 105.695 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.53 0 17.53 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.805 0 72.805 4 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.26 156.505 51.26 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.805 156.505 72.805 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.72 156.505 83.72 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.695 156.505 105.695 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.615 156.505 116.615 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.56 156.505 138.56 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.46 156.505 5.46 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.765 156.505 150.765 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.53 156.505 17.53 160.505 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.76 156.505 28.76 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.46 0 5.46 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.805 0 72.805 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.53 0 17.53 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.72 0 83.72 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.695 0 105.695 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.615 0 116.615 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.765 0 150.765 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.56 0 138.56 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.26 0 51.26 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.76 0 28.76 4 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.26 156.505 51.26 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.805 156.505 72.805 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.72 156.505 83.72 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.695 156.505 105.695 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.615 156.505 116.615 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.56 156.505 138.56 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.76 156.505 28.76 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.765 156.505 150.765 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.53 156.505 17.53 160.505 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.46 156.505 5.46 160.505 ;
    END
  END VDD

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.615 0 26.775 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.615 0 26.775 0.16 ;
    END
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 131.235 0 131.395 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.235 0 131.395 0.16 ;
    END
  END OEB1

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 51.905 0 52.065 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.905 0 52.065 0.16 ;
    END
  END O2[9]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.29 0 52.45 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.29 0 52.45 0.16 ;
    END
  END O2[8]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 36.965 0 37.125 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.965 0 37.125 0.16 ;
    END
  END O2[7]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 37.505 0 37.665 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.505 0 37.665 0.16 ;
    END
  END O2[6]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 37.84 0 38 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.84 0 38 0.16 ;
    END
  END O2[5]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 38.195 0 38.355 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.195 0 38.355 0.16 ;
    END
  END O2[4]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 22.855 0 23.015 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.855 0 23.015 0.16 ;
    END
  END O2[3]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 23.29 0 23.45 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.29 0 23.45 0.16 ;
    END
  END O2[2]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 23.625 0 23.785 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.625 0 23.785 0.16 ;
    END
  END O2[1]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.13 0 65.29 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.13 0 65.29 0.16 ;
    END
  END O2[15]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.48 0 65.64 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.48 0 65.64 0.16 ;
    END
  END O2[14]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.84 0 66 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.84 0 66 0.16 ;
    END
  END O2[13]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.295 0 66.455 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.295 0 66.455 0.16 ;
    END
  END O2[12]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.995 0 51.155 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.995 0 51.155 0.16 ;
    END
  END O2[11]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 51.48 0 51.64 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.48 0 51.64 0.16 ;
    END
  END O2[10]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 23.955 0 24.115 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.955 0 24.115 0.16 ;
    END
  END O2[0]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.01 0 120.17 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.01 0 120.17 0.16 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.655 0 119.815 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 119.655 0 119.815 0.16 ;
    END
  END O1[8]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.855 0 107.015 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.855 0 107.015 0.16 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.37 0 106.53 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.37 0 106.53 0.16 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.945 0 106.105 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.945 0 106.105 0.16 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.56 0 105.72 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.56 0 105.72 0.16 ;
    END
  END O1[4]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.72 0 92.88 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.72 0 92.88 0.16 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.37 0 92.53 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.37 0 92.53 0.16 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.01 0 92.17 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.01 0 92.17 0.16 ;
    END
  END O1[1]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 134.995 0 135.155 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 134.995 0 135.155 0.16 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 134.56 0 134.72 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 134.56 0 134.72 0.16 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 134.225 0 134.385 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 134.225 0 134.385 0.16 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.895 0 134.055 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 133.895 0 134.055 0.16 ;
    END
  END O1[12]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.885 0 121.045 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.885 0 121.045 0.16 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.345 0 120.505 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.345 0 120.505 0.16 ;
    END
  END O1[10]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 91.555 0 91.715 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.555 0 91.715 0.16 ;
    END
  END O1[0]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 56.655 0 56.815 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.655 0 56.815 0.16 ;
    END
  END I2[9]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 56.335 0 56.495 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.335 0 56.495 0.16 ;
    END
  END I2[8]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 43.505 0 43.665 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.505 0 43.665 0.16 ;
    END
  END I2[7]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.895 0 43.055 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.895 0 43.055 0.16 ;
    END
  END I2[6]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.575 0 42.735 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.575 0 42.735 0.16 ;
    END
  END I2[5]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.255 0 42.415 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.255 0 42.415 0.16 ;
    END
  END I2[4]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.425 0 29.585 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.425 0 29.585 0.16 ;
    END
  END I2[3]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.815 0 28.975 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.815 0 28.975 0.16 ;
    END
  END I2[2]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.495 0 28.655 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.495 0 28.655 0.16 ;
    END
  END I2[1]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.665 0 71.825 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.665 0 71.825 0.16 ;
    END
  END I2[15]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.055 0 71.215 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.055 0 71.215 0.16 ;
    END
  END I2[14]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 70.735 0 70.895 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.735 0 70.895 0.16 ;
    END
  END I2[13]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 70.415 0 70.575 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.415 0 70.575 0.16 ;
    END
  END I2[12]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.585 0 57.745 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.585 0 57.745 0.16 ;
    END
  END I2[11]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 56.975 0 57.135 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.975 0 57.135 0.16 ;
    END
  END I2[10]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.175 0 28.335 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.175 0 28.335 0.16 ;
    END
  END I2[0]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.275 0 115.435 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 115.275 0 115.435 0.16 ;
    END
  END I1[9]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.595 0 115.755 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 115.595 0 115.755 0.16 ;
    END
  END I1[8]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.265 0 100.425 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.265 0 100.425 0.16 ;
    END
  END I1[7]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.875 0 101.035 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.875 0 101.035 0.16 ;
    END
  END I1[6]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.195 0 101.355 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.195 0 101.355 0.16 ;
    END
  END I1[5]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.515 0 101.675 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.515 0 101.675 0.16 ;
    END
  END I1[4]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 86.185 0 86.345 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.185 0 86.345 0.16 ;
    END
  END I1[3]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 86.795 0 86.955 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.795 0 86.955 0.16 ;
    END
  END I1[2]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.115 0 87.275 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.115 0 87.275 0.16 ;
    END
  END I1[1]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 128.425 0 128.585 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 128.425 0 128.585 0.16 ;
    END
  END I1[15]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.035 0 129.195 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 129.035 0 129.195 0.16 ;
    END
  END I1[14]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.355 0 129.515 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 129.355 0 129.515 0.16 ;
    END
  END I1[13]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.675 0 129.835 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 129.675 0 129.835 0.16 ;
    END
  END I1[12]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.345 0 114.505 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 114.345 0 114.505 0.16 ;
    END
  END I1[11]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.955 0 115.115 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 114.955 0 115.115 0.16 ;
    END
  END I1[10]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.435 0 87.595 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.435 0 87.595 0.16 ;
    END
  END I1[0]

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 21.93 0 22.09 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.93 0 22.09 0.16 ;
    END
  END CSB2

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.92 0 136.08 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 135.92 0 136.08 0.16 ;
    END
  END CSB1

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 19.33 0 19.49 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 19.33 0 19.49 0.16 ;
    END
  END CE2

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.52 0 138.68 0.16 ;
    END
    PORT
      LAYER M2 ;
        RECT 138.52 0 138.68 0.16 ;
    END
  END CE1

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 96.735 0.16 96.895 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 96.735 0.16 96.895 ;
    END
  END A2[5]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 99.96 0.16 100.12 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 99.96 0.16 100.12 ;
    END
  END A2[4]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 102.54 0.16 102.7 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 102.54 0.16 102.7 ;
    END
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 105.755 0.16 105.915 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 105.755 0.16 105.915 ;
    END
  END A2[2]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 108.255 0.16 108.415 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 108.255 0.16 108.415 ;
    END
  END A2[1]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 111.46 0.275 111.735 ;
    END
    PORT
      LAYER M2 ;
        RECT 0 111.46 0.275 111.735 ;
    END
  END A2[0]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.43 96.75 154.59 96.91 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.43 96.75 154.59 96.91 ;
    END
  END A1[5]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.43 99.96 154.59 100.12 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.43 99.96 154.59 100.12 ;
    END
  END A1[4]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.43 102.54 154.59 102.7 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.43 102.54 154.59 102.7 ;
    END
  END A1[3]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.43 105.755 154.59 105.915 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.43 105.755 154.59 105.915 ;
    END
  END A1[2]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.43 108.255 154.59 108.415 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.43 108.255 154.59 108.415 ;
    END
  END A1[1]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.315 111.46 154.59 111.735 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.315 111.46 154.59 111.735 ;
    END
  END A1[0]
  OBS
    LAYER M3 ;
      RECT 0.32 96.59 154.27 97.055 ;
      RECT 0 111.895 154.59 160.505 ;
      RECT 0 108.575 154.59 111.3 ;
      RECT 0 106.075 154.59 108.095 ;
      RECT 0 102.86 154.59 105.595 ;
      RECT 0 100.28 154.59 102.38 ;
      RECT 0 97.07 154.59 99.8 ;
      RECT 0 35.455 154.59 96.575 ;
      RECT 0 34.385 154.59 34.975 ;
      RECT 0 0.32 154.59 33.905 ;
      RECT 0.435 111.3 154.155 111.895 ;
      RECT 0.32 108.095 154.27 108.575 ;
      RECT 0.32 105.595 154.27 106.075 ;
      RECT 0.32 102.38 154.27 102.86 ;
      RECT 0 97.055 154.27 97.07 ;
      RECT 0.32 99.8 154.27 100.28 ;
      RECT 0.32 96.575 154.59 96.59 ;
      RECT 0.32 34.975 154.59 35.455 ;
      RECT 71.985 0 86.025 0.32 ;
      RECT 138.84 0 154.59 0.32 ;
      RECT 136.24 0 138.36 0.32 ;
      RECT 135.315 0 135.76 0.32 ;
      RECT 129.995 0 131.075 0.32 ;
      RECT 131.555 0 133.735 0.32 ;
      RECT 121.205 0 128.265 0.32 ;
      RECT 115.915 0 119.495 0.32 ;
      RECT 107.175 0 114.185 0.32 ;
      RECT 101.835 0 105.4 0.32 ;
      RECT 93.04 0 100.105 0.32 ;
      RECT 87.755 0 91.395 0.32 ;
      RECT 66.615 0 70.255 0.32 ;
      RECT 57.905 0 64.97 0.32 ;
      RECT 52.61 0 56.175 0.32 ;
      RECT 43.825 0 50.835 0.32 ;
      RECT 38.515 0 42.095 0.32 ;
      RECT 29.745 0 36.805 0.32 ;
      RECT 24.275 0 26.455 0.32 ;
      RECT 26.935 0 28.015 0.32 ;
      RECT 22.25 0 22.695 0.32 ;
      RECT 19.65 0 21.77 0.32 ;
      RECT 0 0 19.17 0.32 ;
      RECT 0 33.905 154.27 34.385 ;
    LAYER M2 ;
      RECT 0 111.895 154.59 160.505 ;
      RECT 0 108.575 154.59 111.3 ;
      RECT 0 106.075 154.59 108.095 ;
      RECT 0 102.86 154.59 105.595 ;
      RECT 0 100.28 154.59 102.38 ;
      RECT 0 97.07 154.59 99.8 ;
      RECT 0 35.455 154.59 96.575 ;
      RECT 0 34.385 154.59 34.975 ;
      RECT 0 0.32 154.59 33.905 ;
      RECT 0.435 111.3 154.155 111.895 ;
      RECT 0.32 108.095 154.27 108.575 ;
      RECT 0.32 105.595 154.27 106.075 ;
      RECT 0.32 102.38 154.27 102.86 ;
      RECT 0 97.055 154.27 97.07 ;
      RECT 0.32 99.8 154.27 100.28 ;
      RECT 0.32 96.575 154.59 96.59 ;
      RECT 0.32 34.975 154.59 35.455 ;
      RECT 71.985 0 86.025 0.32 ;
      RECT 138.84 0 154.59 0.32 ;
      RECT 136.24 0 138.36 0.32 ;
      RECT 135.315 0 135.76 0.32 ;
      RECT 129.995 0 131.075 0.32 ;
      RECT 131.555 0 133.735 0.32 ;
      RECT 121.205 0 128.265 0.32 ;
      RECT 115.915 0 119.495 0.32 ;
      RECT 107.175 0 114.185 0.32 ;
      RECT 101.835 0 105.4 0.32 ;
      RECT 93.04 0 100.105 0.32 ;
      RECT 87.755 0 91.395 0.32 ;
      RECT 66.615 0 70.255 0.32 ;
      RECT 57.905 0 64.97 0.32 ;
      RECT 52.61 0 56.175 0.32 ;
      RECT 43.825 0 50.835 0.32 ;
      RECT 38.515 0 42.095 0.32 ;
      RECT 29.745 0 36.805 0.32 ;
      RECT 24.275 0 26.455 0.32 ;
      RECT 26.935 0 28.015 0.32 ;
      RECT 22.25 0 22.695 0.32 ;
      RECT 19.65 0 21.77 0.32 ;
      RECT 0 0 19.17 0.32 ;
      RECT 0 33.905 154.27 34.385 ;
      RECT 0.32 96.59 154.27 97.055 ;
    LAYER M1 ;
      RECT 0 0 154.59 160.505 ;
    LAYER PO ;
      RECT 0 0 154.59 160.505 ;
    LAYER M5 ;
      RECT 0 4.16 154.59 156.345 ;
      RECT 150.925 156.345 154.59 160.505 ;
      RECT 138.72 156.345 141.295 160.505 ;
      RECT 145.615 156.345 146.605 160.505 ;
      RECT 116.775 156.345 129.09 160.505 ;
      RECT 133.41 156.345 134.4 160.505 ;
      RECT 150.925 0 154.59 4.16 ;
      RECT 138.72 0 141.295 4.16 ;
      RECT 145.615 0 146.605 4.16 ;
      RECT 116.775 0 129.09 4.16 ;
      RECT 133.41 0 134.4 4.16 ;
      RECT 105.855 156.345 107.145 160.505 ;
      RECT 111.465 156.345 112.455 160.505 ;
      RECT 83.88 156.345 96.225 160.505 ;
      RECT 100.545 156.345 101.535 160.505 ;
      RECT 78.57 156.345 79.56 160.505 ;
      RECT 105.855 0 107.145 4.16 ;
      RECT 111.465 0 112.455 4.16 ;
      RECT 83.88 0 96.225 4.16 ;
      RECT 100.545 0 101.535 4.16 ;
      RECT 78.57 0 79.56 4.16 ;
      RECT 28.92 156.345 41.79 160.505 ;
      RECT 28.92 0 41.79 4.16 ;
      RECT 72.965 156.345 74.25 160.505 ;
      RECT 51.42 156.345 63.335 160.505 ;
      RECT 67.655 156.345 68.645 160.505 ;
      RECT 46.11 156.345 47.1 160.505 ;
      RECT 72.965 0 74.25 4.16 ;
      RECT 51.42 0 63.335 4.16 ;
      RECT 67.655 0 68.645 4.16 ;
      RECT 46.11 0 47.1 4.16 ;
      RECT 17.69 156.345 19.29 160.505 ;
      RECT 23.61 156.345 24.6 160.505 ;
      RECT 5.62 156.345 7.25 160.505 ;
      RECT 11.57 156.345 13.37 160.505 ;
      RECT 0 156.345 1.3 160.505 ;
      RECT 17.69 0 19.29 4.16 ;
      RECT 23.61 0 24.6 4.16 ;
      RECT 5.62 0 7.25 4.16 ;
      RECT 11.57 0 13.37 4.16 ;
      RECT 0 0 1.3 4.16 ;
    LAYER M4 ;
      RECT 0 4.16 154.59 156.345 ;
      RECT 150.925 156.345 154.59 160.505 ;
      RECT 138.72 156.345 141.295 160.505 ;
      RECT 145.615 156.345 146.605 160.505 ;
      RECT 116.775 156.345 129.09 160.505 ;
      RECT 133.41 156.345 134.4 160.505 ;
      RECT 150.925 0 154.59 4.16 ;
      RECT 138.72 0 141.295 4.16 ;
      RECT 145.615 0 146.605 4.16 ;
      RECT 116.775 0 129.09 4.16 ;
      RECT 133.41 0 134.4 4.16 ;
      RECT 105.855 156.345 107.145 160.505 ;
      RECT 111.465 156.345 112.455 160.505 ;
      RECT 83.88 156.345 96.225 160.505 ;
      RECT 100.545 156.345 101.535 160.505 ;
      RECT 78.57 156.345 79.56 160.505 ;
      RECT 105.855 0 107.145 4.16 ;
      RECT 111.465 0 112.455 4.16 ;
      RECT 83.88 0 96.225 4.16 ;
      RECT 100.545 0 101.535 4.16 ;
      RECT 78.57 0 79.56 4.16 ;
      RECT 28.92 156.345 41.79 160.505 ;
      RECT 28.92 0 41.79 4.16 ;
      RECT 72.965 156.345 74.25 160.505 ;
      RECT 51.42 156.345 63.335 160.505 ;
      RECT 67.655 156.345 68.645 160.505 ;
      RECT 46.11 156.345 47.1 160.505 ;
      RECT 72.965 0 74.25 4.16 ;
      RECT 51.42 0 63.335 4.16 ;
      RECT 67.655 0 68.645 4.16 ;
      RECT 46.11 0 47.1 4.16 ;
      RECT 17.69 156.345 19.29 160.505 ;
      RECT 23.61 156.345 24.6 160.505 ;
      RECT 5.62 156.345 7.25 160.505 ;
      RECT 11.57 156.345 13.37 160.505 ;
      RECT 0 156.345 1.3 160.505 ;
      RECT 17.69 0 19.29 4.16 ;
      RECT 23.61 0 24.6 4.16 ;
      RECT 5.62 0 7.25 4.16 ;
      RECT 11.57 0 13.37 4.16 ;
      RECT 0 0 1.3 4.16 ;
  END
END SRAM16x64
  
END LIBRARY
